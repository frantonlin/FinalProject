`timescale 1 ns / 1 ps
`include "fpuAdder.v"

module testFpuAdder();
    wire [31:0] Z;
    reg op;
    reg [31:0] A, B;

    fpuAdder fpuAdder0(Z, op, A, B);

    initial begin
        $dumpfile("fpuAdder_all.vcd");
        $dumpvars();

        $display("A                     op    B                    =  Z");
        A=32'b01000000000000000000000000000000;
        B=32'b01000000010000000000000000000000;
        op=0;#1000;
        $display("%s * 2^%-1d * %f  %s  %s * 2^%-1d * %f  =  %s * 2^%-1d * %f    %b", A[31]?"-1":"+1",$signed(A[30:23]-127),$itor({1'b1,A[22:0]})*(2.0**-23.0), op?"MINUS":"PLUS", B[31]?"-1":"+1",$signed(B[30:23]-127),$itor({1'b1,B[22:0]})*(2.0**-23.0), Z[31]?"-1":"+1",$signed(Z[30:23]-127),$itor({1'b1,Z[22:0]})*(2.0**-23.0), Z);
        $display("%f %s %f = %f", $itor((A[31]?-1:1)*2**(A[30:23]-127)*{1'b1,A[22:0]})*(2.0**-23.0),  op?"-":"+", $itor((B[31]?-1:1)*2**(B[30:23]-127)*{1'b1,B[22:0]})*(2.0**-23.0), $itor((Z[31]?-1:1)*2**(Z[30:23]-127)*{1'b1,Z[22:0]})*(2.0**-23.0));
        $display();

        A=32'b11000000000000000000000000000000;
        B=32'b11000000010000000000000000000000;
        op=1;#1000;
        $display("%s * 2^%-1d * %f  %s  %s * 2^%-1d * %f  =  %s * 2^%-1d * %f    %b", A[31]?"-1":"+1",$signed(A[30:23]-127),$itor({1'b1,A[22:0]})*(2.0**-23.0), op?"MINUS":"PLUS", B[31]?"-1":"+1",$signed(B[30:23]-127),$itor({1'b1,B[22:0]})*(2.0**-23.0), Z[31]?"-1":"+1",$signed(Z[30:23]-127),$itor({1'b1,Z[22:0]})*(2.0**-23.0), Z);
        $display("%f %s %f = %f", $itor((A[31]?-1:1)*2**(A[30:23]-127)*{1'b1,A[22:0]})*(2.0**-23.0),  op?"-":"+", $itor((B[31]?-1:1)*2**(B[30:23]-127)*{1'b1,B[22:0]})*(2.0**-23.0), $itor((Z[31]?-1:1)*2**(Z[30:23]-127)*{1'b1,Z[22:0]})*(2.0**-23.0));
        $display();

        A=32'b00111111000000000000000000000000; //0.5
        B=32'b00111111000000000000000000000000; //0.5
        op=0;#1000;
        $display("%s * 2^%-1d * %f  %s  %s * 2^%-1d * %f  =  %s * 2^%-1d * %f    %b", A[31]?"-1":"+1",$signed(A[30:23]-127),$itor({1'b1,A[22:0]})*(2.0**-23.0), op?"MINUS":"PLUS", B[31]?"-1":"+1",$signed(B[30:23]-127),$itor({1'b1,B[22:0]})*(2.0**-23.0), Z[31]?"-1":"+1",$signed(Z[30:23]-127),$itor({1'b1,Z[22:0]})*(2.0**-23.0), Z);
        $display("%f %s %f = %f", (A[31]?-1:1)*2**(A[30:23]-127)*{1'b1,A[22:0]}*(2.0**-23.0),  op?"-":"+", $itor((B[31]?-1:1)*2**(B[30:23]-127)*{1'b1,B[22:0]})*(2.0**-23.0), $itor((Z[31]?-1:1)*2**(Z[30:23]-127)*{1'b1,Z[22:0]})*(2.0**-23.0));

        $dumpflush;
    end

endmodule

